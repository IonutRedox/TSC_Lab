/***********************************************************************
 * A SystemVerilog RTL model of an instruction register:
 * User-defined type definitions
 **********************************************************************/
package instr_register_test_pkg;
  `include "driver.sv";
  `include "transaction.sv";
  `include "monitor.sv";
endpackage
